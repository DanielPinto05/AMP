package 
    parameter logic[3:0] OP_ADD = 4'b0000;
    parameter logic[3:0] OP_SUB = 4'b0001;
    parameter logic[3:0] OP_SLL = 4'b0010;
    parameter logic[3:0] OP_SRA = 4'b0011;
    parameter logic[3:0] OP_SRL = 4'b0100;
    parameter logic[3:0] OP_OR = 4'b0101;
    parameter logic[3:0] OP_XOR = 4'b0110;
    parameter logic[3:0] OP_SSLT = 4'b0111;
    parameter logic[3:0] OP_USLT = 4'b1000;
    parameter logic[3:0] OP_AND = 4'b1001;
    
endpackage