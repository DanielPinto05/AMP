module FSM(
    input logic op[6:0], 
    input logic funct7_5; 
    input logic funct3[2:0]; 
);

endmodule